module GunControl();

endmodule 

module test (
	clk_clk,
	reset_reset_n,
	led_pio_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	led_pio_external_connection_export;
endmodule

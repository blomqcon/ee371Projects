library verilog;
use verilog.vl_types.all;
entity mux4_1_testbench is
end mux4_1_testbench;

module GameTime();

endmodule
module AliensControl();

endmodule 
module BitIdentifierCount(identifer, enable, bscClk);
	input enable, bscClk;
	output [7:0] identifer;
	
endmodule 
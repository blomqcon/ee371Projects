library verilog;
use verilog.vl_types.all;
entity DE1_SoC_testbench is
end DE1_SoC_testbench;

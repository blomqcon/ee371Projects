// nios_system.v

// Generated using ACDS version 14.0 200 at 2016.03.04.18:44:50

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        reset_reset_n,                                               //                                                reset.reset_n
		input  wire [7:0]  receive_parallel_to_processor_external_connection_export,    //    receive_parallel_to_processor_external_connection.export
		input  wire        clk_clk,                                                     //                                                  clk.clk
		output wire [7:0]  transmit_parallel_from_processor_external_connection_export, // transmit_parallel_from_processor_external_connection.export
		output wire        transmit_enable_external_connection_export,                  //                  transmit_enable_external_connection.export
		input  wire        transmit_character_sent_external_connection_export,          //          transmit_character_sent_external_connection.export
		output wire        transmit_load_external_connection_export,                    //                    transmit_load_external_connection.export
		input  wire        received_character_received_external_connection_export,      //      received_character_received_external_connection.export
		output wire [10:0] sram_address_external_connection_export,                     //                     sram_address_external_connection.export
		inout  wire [7:0]  sram_data_external_connection_export,                        //                        sram_data_external_connection.export
		output wire        sram_enable_external_connection_export,                      //                      sram_enable_external_connection.export
		output wire        sram_read_write_external_connection_export,                  //                  sram_read_write_external_connection.export
		input  wire        gunner_left_external_connection_export,                      //                      gunner_left_external_connection.export
		input  wire        gunner_right_external_connection_export,                     //                     gunner_right_external_connection.export
		input  wire [1:0]  gunner_shoot_external_connection_export,                     //                     gunner_shoot_external_connection.export
		input  wire        alien_shoot_external_connection_export,                      //                      alien_shoot_external_connection.export
		input  wire [2:0]  alien_x_position_external_connection_export,                 //                 alien_x_position_external_connection.export
		input  wire [1:0]  alien_y_position_external_connection_export,                 //                 alien_y_position_external_connection.export
		input  wire [31:0] game_timer_external_connection_export,                       //                       game_timer_external_connection.export
		input  wire [15:0] random_number_lfsr_output_external_connection_export         //        random_number_lfsr_output_external_connection.export
	);

	wire         cpu_instruction_master_waitrequest;                               // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [13:0] cpu_instruction_master_address;                                   // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                      // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                  // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_data_master_waitrequest;                                      // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                        // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [13:0] cpu_data_master_address;                                          // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                            // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                             // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                         // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                      // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                       // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;              // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                  // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                    // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                     // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                 // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;              // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;               // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;                    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                 // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                 // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;      // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;            // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;             // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;         // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire   [1:0] mm_interconnect_0_receive_parallel_to_processor_s1_address;       // mm_interconnect_0:RECEIVE_PARALLEL_TO_PROCESSOR_s1_address -> RECEIVE_PARALLEL_TO_PROCESSOR:address
	wire  [31:0] mm_interconnect_0_receive_parallel_to_processor_s1_readdata;      // RECEIVE_PARALLEL_TO_PROCESSOR:readdata -> mm_interconnect_0:RECEIVE_PARALLEL_TO_PROCESSOR_s1_readdata
	wire  [31:0] mm_interconnect_0_transmit_parallel_from_processor_s1_writedata;  // mm_interconnect_0:TRANSMIT_PARALLEL_FROM_PROCESSOR_s1_writedata -> TRANSMIT_PARALLEL_FROM_PROCESSOR:writedata
	wire   [1:0] mm_interconnect_0_transmit_parallel_from_processor_s1_address;    // mm_interconnect_0:TRANSMIT_PARALLEL_FROM_PROCESSOR_s1_address -> TRANSMIT_PARALLEL_FROM_PROCESSOR:address
	wire         mm_interconnect_0_transmit_parallel_from_processor_s1_chipselect; // mm_interconnect_0:TRANSMIT_PARALLEL_FROM_PROCESSOR_s1_chipselect -> TRANSMIT_PARALLEL_FROM_PROCESSOR:chipselect
	wire         mm_interconnect_0_transmit_parallel_from_processor_s1_write;      // mm_interconnect_0:TRANSMIT_PARALLEL_FROM_PROCESSOR_s1_write -> TRANSMIT_PARALLEL_FROM_PROCESSOR:write_n
	wire  [31:0] mm_interconnect_0_transmit_parallel_from_processor_s1_readdata;   // TRANSMIT_PARALLEL_FROM_PROCESSOR:readdata -> mm_interconnect_0:TRANSMIT_PARALLEL_FROM_PROCESSOR_s1_readdata
	wire  [31:0] mm_interconnect_0_transmit_enable_s1_writedata;                   // mm_interconnect_0:TRANSMIT_ENABLE_s1_writedata -> TRANSMIT_ENABLE:writedata
	wire   [1:0] mm_interconnect_0_transmit_enable_s1_address;                     // mm_interconnect_0:TRANSMIT_ENABLE_s1_address -> TRANSMIT_ENABLE:address
	wire         mm_interconnect_0_transmit_enable_s1_chipselect;                  // mm_interconnect_0:TRANSMIT_ENABLE_s1_chipselect -> TRANSMIT_ENABLE:chipselect
	wire         mm_interconnect_0_transmit_enable_s1_write;                       // mm_interconnect_0:TRANSMIT_ENABLE_s1_write -> TRANSMIT_ENABLE:write_n
	wire  [31:0] mm_interconnect_0_transmit_enable_s1_readdata;                    // TRANSMIT_ENABLE:readdata -> mm_interconnect_0:TRANSMIT_ENABLE_s1_readdata
	wire   [1:0] mm_interconnect_0_transmit_character_sent_s1_address;             // mm_interconnect_0:TRANSMIT_CHARACTER_SENT_s1_address -> TRANSMIT_CHARACTER_SENT:address
	wire  [31:0] mm_interconnect_0_transmit_character_sent_s1_readdata;            // TRANSMIT_CHARACTER_SENT:readdata -> mm_interconnect_0:TRANSMIT_CHARACTER_SENT_s1_readdata
	wire  [31:0] mm_interconnect_0_transmit_load_s1_writedata;                     // mm_interconnect_0:TRANSMIT_LOAD_s1_writedata -> TRANSMIT_LOAD:writedata
	wire   [1:0] mm_interconnect_0_transmit_load_s1_address;                       // mm_interconnect_0:TRANSMIT_LOAD_s1_address -> TRANSMIT_LOAD:address
	wire         mm_interconnect_0_transmit_load_s1_chipselect;                    // mm_interconnect_0:TRANSMIT_LOAD_s1_chipselect -> TRANSMIT_LOAD:chipselect
	wire         mm_interconnect_0_transmit_load_s1_write;                         // mm_interconnect_0:TRANSMIT_LOAD_s1_write -> TRANSMIT_LOAD:write_n
	wire  [31:0] mm_interconnect_0_transmit_load_s1_readdata;                      // TRANSMIT_LOAD:readdata -> mm_interconnect_0:TRANSMIT_LOAD_s1_readdata
	wire   [1:0] mm_interconnect_0_receive_character_received_s1_address;          // mm_interconnect_0:RECEIVE_CHARACTER_RECEIVED_s1_address -> RECEIVE_CHARACTER_RECEIVED:address
	wire  [31:0] mm_interconnect_0_receive_character_received_s1_readdata;         // RECEIVE_CHARACTER_RECEIVED:readdata -> mm_interconnect_0:RECEIVE_CHARACTER_RECEIVED_s1_readdata
	wire  [31:0] mm_interconnect_0_sram_address_s1_writedata;                      // mm_interconnect_0:SRAM_ADDRESS_s1_writedata -> SRAM_ADDRESS:writedata
	wire   [1:0] mm_interconnect_0_sram_address_s1_address;                        // mm_interconnect_0:SRAM_ADDRESS_s1_address -> SRAM_ADDRESS:address
	wire         mm_interconnect_0_sram_address_s1_chipselect;                     // mm_interconnect_0:SRAM_ADDRESS_s1_chipselect -> SRAM_ADDRESS:chipselect
	wire         mm_interconnect_0_sram_address_s1_write;                          // mm_interconnect_0:SRAM_ADDRESS_s1_write -> SRAM_ADDRESS:write_n
	wire  [31:0] mm_interconnect_0_sram_address_s1_readdata;                       // SRAM_ADDRESS:readdata -> mm_interconnect_0:SRAM_ADDRESS_s1_readdata
	wire  [31:0] mm_interconnect_0_sram_data_s1_writedata;                         // mm_interconnect_0:SRAM_DATA_s1_writedata -> SRAM_DATA:writedata
	wire   [1:0] mm_interconnect_0_sram_data_s1_address;                           // mm_interconnect_0:SRAM_DATA_s1_address -> SRAM_DATA:address
	wire         mm_interconnect_0_sram_data_s1_chipselect;                        // mm_interconnect_0:SRAM_DATA_s1_chipselect -> SRAM_DATA:chipselect
	wire         mm_interconnect_0_sram_data_s1_write;                             // mm_interconnect_0:SRAM_DATA_s1_write -> SRAM_DATA:write_n
	wire  [31:0] mm_interconnect_0_sram_data_s1_readdata;                          // SRAM_DATA:readdata -> mm_interconnect_0:SRAM_DATA_s1_readdata
	wire  [31:0] mm_interconnect_0_sram_enable_s1_writedata;                       // mm_interconnect_0:SRAM_ENABLE_s1_writedata -> SRAM_ENABLE:writedata
	wire   [1:0] mm_interconnect_0_sram_enable_s1_address;                         // mm_interconnect_0:SRAM_ENABLE_s1_address -> SRAM_ENABLE:address
	wire         mm_interconnect_0_sram_enable_s1_chipselect;                      // mm_interconnect_0:SRAM_ENABLE_s1_chipselect -> SRAM_ENABLE:chipselect
	wire         mm_interconnect_0_sram_enable_s1_write;                           // mm_interconnect_0:SRAM_ENABLE_s1_write -> SRAM_ENABLE:write_n
	wire  [31:0] mm_interconnect_0_sram_enable_s1_readdata;                        // SRAM_ENABLE:readdata -> mm_interconnect_0:SRAM_ENABLE_s1_readdata
	wire  [31:0] mm_interconnect_0_sram_read_write_s1_writedata;                   // mm_interconnect_0:SRAM_READ_WRITE_s1_writedata -> SRAM_READ_WRITE:writedata
	wire   [1:0] mm_interconnect_0_sram_read_write_s1_address;                     // mm_interconnect_0:SRAM_READ_WRITE_s1_address -> SRAM_READ_WRITE:address
	wire         mm_interconnect_0_sram_read_write_s1_chipselect;                  // mm_interconnect_0:SRAM_READ_WRITE_s1_chipselect -> SRAM_READ_WRITE:chipselect
	wire         mm_interconnect_0_sram_read_write_s1_write;                       // mm_interconnect_0:SRAM_READ_WRITE_s1_write -> SRAM_READ_WRITE:write_n
	wire  [31:0] mm_interconnect_0_sram_read_write_s1_readdata;                    // SRAM_READ_WRITE:readdata -> mm_interconnect_0:SRAM_READ_WRITE_s1_readdata
	wire   [1:0] mm_interconnect_0_gunner_left_s1_address;                         // mm_interconnect_0:GUNNER_LEFT_s1_address -> GUNNER_LEFT:address
	wire  [31:0] mm_interconnect_0_gunner_left_s1_readdata;                        // GUNNER_LEFT:readdata -> mm_interconnect_0:GUNNER_LEFT_s1_readdata
	wire   [1:0] mm_interconnect_0_gunner_right_s1_address;                        // mm_interconnect_0:GUNNER_RIGHT_s1_address -> GUNNER_RIGHT:address
	wire  [31:0] mm_interconnect_0_gunner_right_s1_readdata;                       // GUNNER_RIGHT:readdata -> mm_interconnect_0:GUNNER_RIGHT_s1_readdata
	wire   [1:0] mm_interconnect_0_gunner_shoot_s1_address;                        // mm_interconnect_0:GUNNER_SHOOT_s1_address -> GUNNER_SHOOT:address
	wire  [31:0] mm_interconnect_0_gunner_shoot_s1_readdata;                       // GUNNER_SHOOT:readdata -> mm_interconnect_0:GUNNER_SHOOT_s1_readdata
	wire   [1:0] mm_interconnect_0_alien_shoot_s1_address;                         // mm_interconnect_0:ALIEN_SHOOT_s1_address -> ALIEN_SHOOT:address
	wire  [31:0] mm_interconnect_0_alien_shoot_s1_readdata;                        // ALIEN_SHOOT:readdata -> mm_interconnect_0:ALIEN_SHOOT_s1_readdata
	wire   [1:0] mm_interconnect_0_alien_x_position_s1_address;                    // mm_interconnect_0:ALIEN_X_POSITION_s1_address -> ALIEN_X_POSITION:address
	wire  [31:0] mm_interconnect_0_alien_x_position_s1_readdata;                   // ALIEN_X_POSITION:readdata -> mm_interconnect_0:ALIEN_X_POSITION_s1_readdata
	wire   [1:0] mm_interconnect_0_alien_y_position_s1_address;                    // mm_interconnect_0:ALIEN_Y_POSITION_s1_address -> ALIEN_Y_POSITION:address
	wire  [31:0] mm_interconnect_0_alien_y_position_s1_readdata;                   // ALIEN_Y_POSITION:readdata -> mm_interconnect_0:ALIEN_Y_POSITION_s1_readdata
	wire   [1:0] mm_interconnect_0_game_timer_s1_address;                          // mm_interconnect_0:GAME_TIMER_s1_address -> GAME_TIMER:address
	wire  [31:0] mm_interconnect_0_game_timer_s1_readdata;                         // GAME_TIMER:readdata -> mm_interconnect_0:GAME_TIMER_s1_readdata
	wire   [1:0] mm_interconnect_0_random_number_lfsr_output_s1_address;           // mm_interconnect_0:RANDOM_NUMBER_LFSR_OUTPUT_s1_address -> RANDOM_NUMBER_LFSR_OUTPUT:address
	wire  [31:0] mm_interconnect_0_random_number_lfsr_output_s1_readdata;          // RANDOM_NUMBER_LFSR_OUTPUT:readdata -> mm_interconnect_0:RANDOM_NUMBER_LFSR_OUTPUT_s1_readdata
	wire         irq_mapper_receiver0_irq;                                         // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_d_irq_irq;                                                    // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [ALIEN_SHOOT:reset_n, ALIEN_X_POSITION:reset_n, ALIEN_Y_POSITION:reset_n, GAME_TIMER:reset_n, GUNNER_LEFT:reset_n, GUNNER_RIGHT:reset_n, GUNNER_SHOOT:reset_n, RANDOM_NUMBER_LFSR_OUTPUT:reset_n, RECEIVE_CHARACTER_RECEIVED:reset_n, RECEIVE_PARALLEL_TO_PROCESSOR:reset_n, SRAM_ADDRESS:reset_n, SRAM_DATA:reset_n, SRAM_ENABLE:reset_n, SRAM_READ_WRITE:reset_n, TRANSMIT_CHARACTER_SENT:reset_n, TRANSMIT_ENABLE:reset_n, TRANSMIT_LOAD:reset_n, TRANSMIT_PARALLEL_FROM_PROCESSOR:reset_n, cpu:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                               // rst_controller:reset_req -> [cpu:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                                // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	nios_system_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_RECEIVE_PARALLEL_TO_PROCESSOR receive_parallel_to_processor (
		.clk      (clk_clk),                                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                             //               reset.reset_n
		.address  (mm_interconnect_0_receive_parallel_to_processor_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_receive_parallel_to_processor_s1_readdata), //                    .readdata
		.in_port  (receive_parallel_to_processor_external_connection_export)     // external_connection.export
	);

	nios_system_TRANSMIT_PARALLEL_FROM_PROCESSOR transmit_parallel_from_processor (
		.clk        (clk_clk),                                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                                  //               reset.reset_n
		.address    (mm_interconnect_0_transmit_parallel_from_processor_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_transmit_parallel_from_processor_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_transmit_parallel_from_processor_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_transmit_parallel_from_processor_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_transmit_parallel_from_processor_s1_readdata),   //                    .readdata
		.out_port   (transmit_parallel_from_processor_external_connection_export)       // external_connection.export
	);

	nios_system_TRANSMIT_ENABLE transmit_enable (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_transmit_enable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_transmit_enable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_transmit_enable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_transmit_enable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_transmit_enable_s1_readdata),   //                    .readdata
		.out_port   (transmit_enable_external_connection_export)       // external_connection.export
	);

	nios_system_TRANSMIT_CHARACTER_SENT transmit_character_sent (
		.clk      (clk_clk),                                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address  (mm_interconnect_0_transmit_character_sent_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_transmit_character_sent_s1_readdata), //                    .readdata
		.in_port  (transmit_character_sent_external_connection_export)     // external_connection.export
	);

	nios_system_TRANSMIT_ENABLE transmit_load (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_transmit_load_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_transmit_load_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_transmit_load_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_transmit_load_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_transmit_load_s1_readdata),   //                    .readdata
		.out_port   (transmit_load_external_connection_export)       // external_connection.export
	);

	nios_system_TRANSMIT_CHARACTER_SENT receive_character_received (
		.clk      (clk_clk),                                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                          //               reset.reset_n
		.address  (mm_interconnect_0_receive_character_received_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_receive_character_received_s1_readdata), //                    .readdata
		.in_port  (received_character_received_external_connection_export)    // external_connection.export
	);

	nios_system_SRAM_ADDRESS sram_address (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_sram_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sram_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sram_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sram_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sram_address_s1_readdata),   //                    .readdata
		.out_port   (sram_address_external_connection_export)       // external_connection.export
	);

	nios_system_SRAM_DATA sram_data (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_sram_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sram_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sram_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sram_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sram_data_s1_readdata),   //                    .readdata
		.bidir_port (sram_data_external_connection_export)       // external_connection.export
	);

	nios_system_TRANSMIT_ENABLE sram_enable (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_sram_enable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sram_enable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sram_enable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sram_enable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sram_enable_s1_readdata),   //                    .readdata
		.out_port   (sram_enable_external_connection_export)       // external_connection.export
	);

	nios_system_TRANSMIT_ENABLE sram_read_write (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_sram_read_write_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sram_read_write_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sram_read_write_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sram_read_write_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sram_read_write_s1_readdata),   //                    .readdata
		.out_port   (sram_read_write_external_connection_export)       // external_connection.export
	);

	nios_system_TRANSMIT_CHARACTER_SENT gunner_left (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_gunner_left_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_gunner_left_s1_readdata), //                    .readdata
		.in_port  (gunner_left_external_connection_export)     // external_connection.export
	);

	nios_system_TRANSMIT_CHARACTER_SENT gunner_right (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_gunner_right_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_gunner_right_s1_readdata), //                    .readdata
		.in_port  (gunner_right_external_connection_export)     // external_connection.export
	);

	nios_system_GUNNER_SHOOT gunner_shoot (
		.clk      (clk_clk),                                    //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address  (mm_interconnect_0_gunner_shoot_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_gunner_shoot_s1_readdata), //                    .readdata
		.in_port  (gunner_shoot_external_connection_export)     // external_connection.export
	);

	nios_system_TRANSMIT_CHARACTER_SENT alien_shoot (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_alien_shoot_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_alien_shoot_s1_readdata), //                    .readdata
		.in_port  (alien_shoot_external_connection_export)     // external_connection.export
	);

	nios_system_ALIEN_X_POSITION alien_x_position (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_alien_x_position_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_alien_x_position_s1_readdata), //                    .readdata
		.in_port  (alien_x_position_external_connection_export)     // external_connection.export
	);

	nios_system_GUNNER_SHOOT alien_y_position (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_0_alien_y_position_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_alien_y_position_s1_readdata), //                    .readdata
		.in_port  (alien_y_position_external_connection_export)     // external_connection.export
	);

	nios_system_GAME_TIMER game_timer (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_game_timer_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_game_timer_s1_readdata), //                    .readdata
		.in_port  (game_timer_external_connection_export)     // external_connection.export
	);

	nios_system_RANDOM_NUMBER_LFSR_OUTPUT random_number_lfsr_output (
		.clk      (clk_clk),                                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address  (mm_interconnect_0_random_number_lfsr_output_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_random_number_lfsr_output_s1_readdata), //                    .readdata
		.in_port  (random_number_lfsr_output_external_connection_export)     // external_connection.export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                          //                           clk_0_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                                   //   cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                        (cpu_data_master_address),                                          //                     cpu_data_master.address
		.cpu_data_master_waitrequest                    (cpu_data_master_waitrequest),                                      //                                    .waitrequest
		.cpu_data_master_byteenable                     (cpu_data_master_byteenable),                                       //                                    .byteenable
		.cpu_data_master_read                           (cpu_data_master_read),                                             //                                    .read
		.cpu_data_master_readdata                       (cpu_data_master_readdata),                                         //                                    .readdata
		.cpu_data_master_write                          (cpu_data_master_write),                                            //                                    .write
		.cpu_data_master_writedata                      (cpu_data_master_writedata),                                        //                                    .writedata
		.cpu_data_master_debugaccess                    (cpu_data_master_debugaccess),                                      //                                    .debugaccess
		.cpu_instruction_master_address                 (cpu_instruction_master_address),                                   //              cpu_instruction_master.address
		.cpu_instruction_master_waitrequest             (cpu_instruction_master_waitrequest),                               //                                    .waitrequest
		.cpu_instruction_master_read                    (cpu_instruction_master_read),                                      //                                    .read
		.cpu_instruction_master_readdata                (cpu_instruction_master_readdata),                                  //                                    .readdata
		.ALIEN_SHOOT_s1_address                         (mm_interconnect_0_alien_shoot_s1_address),                         //                      ALIEN_SHOOT_s1.address
		.ALIEN_SHOOT_s1_readdata                        (mm_interconnect_0_alien_shoot_s1_readdata),                        //                                    .readdata
		.ALIEN_X_POSITION_s1_address                    (mm_interconnect_0_alien_x_position_s1_address),                    //                 ALIEN_X_POSITION_s1.address
		.ALIEN_X_POSITION_s1_readdata                   (mm_interconnect_0_alien_x_position_s1_readdata),                   //                                    .readdata
		.ALIEN_Y_POSITION_s1_address                    (mm_interconnect_0_alien_y_position_s1_address),                    //                 ALIEN_Y_POSITION_s1.address
		.ALIEN_Y_POSITION_s1_readdata                   (mm_interconnect_0_alien_y_position_s1_readdata),                   //                                    .readdata
		.cpu_jtag_debug_module_address                  (mm_interconnect_0_cpu_jtag_debug_module_address),                  //               cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                    (mm_interconnect_0_cpu_jtag_debug_module_write),                    //                                    .write
		.cpu_jtag_debug_module_read                     (mm_interconnect_0_cpu_jtag_debug_module_read),                     //                                    .read
		.cpu_jtag_debug_module_readdata                 (mm_interconnect_0_cpu_jtag_debug_module_readdata),                 //                                    .readdata
		.cpu_jtag_debug_module_writedata                (mm_interconnect_0_cpu_jtag_debug_module_writedata),                //                                    .writedata
		.cpu_jtag_debug_module_byteenable               (mm_interconnect_0_cpu_jtag_debug_module_byteenable),               //                                    .byteenable
		.cpu_jtag_debug_module_waitrequest              (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),              //                                    .waitrequest
		.cpu_jtag_debug_module_debugaccess              (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),              //                                    .debugaccess
		.GAME_TIMER_s1_address                          (mm_interconnect_0_game_timer_s1_address),                          //                       GAME_TIMER_s1.address
		.GAME_TIMER_s1_readdata                         (mm_interconnect_0_game_timer_s1_readdata),                         //                                    .readdata
		.GUNNER_LEFT_s1_address                         (mm_interconnect_0_gunner_left_s1_address),                         //                      GUNNER_LEFT_s1.address
		.GUNNER_LEFT_s1_readdata                        (mm_interconnect_0_gunner_left_s1_readdata),                        //                                    .readdata
		.GUNNER_RIGHT_s1_address                        (mm_interconnect_0_gunner_right_s1_address),                        //                     GUNNER_RIGHT_s1.address
		.GUNNER_RIGHT_s1_readdata                       (mm_interconnect_0_gunner_right_s1_readdata),                       //                                    .readdata
		.GUNNER_SHOOT_s1_address                        (mm_interconnect_0_gunner_shoot_s1_address),                        //                     GUNNER_SHOOT_s1.address
		.GUNNER_SHOOT_s1_readdata                       (mm_interconnect_0_gunner_shoot_s1_readdata),                       //                                    .readdata
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),          //       jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),            //                                    .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),             //                                    .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),         //                                    .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),        //                                    .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),      //                                    .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),       //                                    .chipselect
		.onchip_memory2_0_s1_address                    (mm_interconnect_0_onchip_memory2_0_s1_address),                    //                 onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                      (mm_interconnect_0_onchip_memory2_0_s1_write),                      //                                    .write
		.onchip_memory2_0_s1_readdata                   (mm_interconnect_0_onchip_memory2_0_s1_readdata),                   //                                    .readdata
		.onchip_memory2_0_s1_writedata                  (mm_interconnect_0_onchip_memory2_0_s1_writedata),                  //                                    .writedata
		.onchip_memory2_0_s1_byteenable                 (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                 //                                    .byteenable
		.onchip_memory2_0_s1_chipselect                 (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                 //                                    .chipselect
		.onchip_memory2_0_s1_clken                      (mm_interconnect_0_onchip_memory2_0_s1_clken),                      //                                    .clken
		.RANDOM_NUMBER_LFSR_OUTPUT_s1_address           (mm_interconnect_0_random_number_lfsr_output_s1_address),           //        RANDOM_NUMBER_LFSR_OUTPUT_s1.address
		.RANDOM_NUMBER_LFSR_OUTPUT_s1_readdata          (mm_interconnect_0_random_number_lfsr_output_s1_readdata),          //                                    .readdata
		.RECEIVE_CHARACTER_RECEIVED_s1_address          (mm_interconnect_0_receive_character_received_s1_address),          //       RECEIVE_CHARACTER_RECEIVED_s1.address
		.RECEIVE_CHARACTER_RECEIVED_s1_readdata         (mm_interconnect_0_receive_character_received_s1_readdata),         //                                    .readdata
		.RECEIVE_PARALLEL_TO_PROCESSOR_s1_address       (mm_interconnect_0_receive_parallel_to_processor_s1_address),       //    RECEIVE_PARALLEL_TO_PROCESSOR_s1.address
		.RECEIVE_PARALLEL_TO_PROCESSOR_s1_readdata      (mm_interconnect_0_receive_parallel_to_processor_s1_readdata),      //                                    .readdata
		.SRAM_ADDRESS_s1_address                        (mm_interconnect_0_sram_address_s1_address),                        //                     SRAM_ADDRESS_s1.address
		.SRAM_ADDRESS_s1_write                          (mm_interconnect_0_sram_address_s1_write),                          //                                    .write
		.SRAM_ADDRESS_s1_readdata                       (mm_interconnect_0_sram_address_s1_readdata),                       //                                    .readdata
		.SRAM_ADDRESS_s1_writedata                      (mm_interconnect_0_sram_address_s1_writedata),                      //                                    .writedata
		.SRAM_ADDRESS_s1_chipselect                     (mm_interconnect_0_sram_address_s1_chipselect),                     //                                    .chipselect
		.SRAM_DATA_s1_address                           (mm_interconnect_0_sram_data_s1_address),                           //                        SRAM_DATA_s1.address
		.SRAM_DATA_s1_write                             (mm_interconnect_0_sram_data_s1_write),                             //                                    .write
		.SRAM_DATA_s1_readdata                          (mm_interconnect_0_sram_data_s1_readdata),                          //                                    .readdata
		.SRAM_DATA_s1_writedata                         (mm_interconnect_0_sram_data_s1_writedata),                         //                                    .writedata
		.SRAM_DATA_s1_chipselect                        (mm_interconnect_0_sram_data_s1_chipselect),                        //                                    .chipselect
		.SRAM_ENABLE_s1_address                         (mm_interconnect_0_sram_enable_s1_address),                         //                      SRAM_ENABLE_s1.address
		.SRAM_ENABLE_s1_write                           (mm_interconnect_0_sram_enable_s1_write),                           //                                    .write
		.SRAM_ENABLE_s1_readdata                        (mm_interconnect_0_sram_enable_s1_readdata),                        //                                    .readdata
		.SRAM_ENABLE_s1_writedata                       (mm_interconnect_0_sram_enable_s1_writedata),                       //                                    .writedata
		.SRAM_ENABLE_s1_chipselect                      (mm_interconnect_0_sram_enable_s1_chipselect),                      //                                    .chipselect
		.SRAM_READ_WRITE_s1_address                     (mm_interconnect_0_sram_read_write_s1_address),                     //                  SRAM_READ_WRITE_s1.address
		.SRAM_READ_WRITE_s1_write                       (mm_interconnect_0_sram_read_write_s1_write),                       //                                    .write
		.SRAM_READ_WRITE_s1_readdata                    (mm_interconnect_0_sram_read_write_s1_readdata),                    //                                    .readdata
		.SRAM_READ_WRITE_s1_writedata                   (mm_interconnect_0_sram_read_write_s1_writedata),                   //                                    .writedata
		.SRAM_READ_WRITE_s1_chipselect                  (mm_interconnect_0_sram_read_write_s1_chipselect),                  //                                    .chipselect
		.TRANSMIT_CHARACTER_SENT_s1_address             (mm_interconnect_0_transmit_character_sent_s1_address),             //          TRANSMIT_CHARACTER_SENT_s1.address
		.TRANSMIT_CHARACTER_SENT_s1_readdata            (mm_interconnect_0_transmit_character_sent_s1_readdata),            //                                    .readdata
		.TRANSMIT_ENABLE_s1_address                     (mm_interconnect_0_transmit_enable_s1_address),                     //                  TRANSMIT_ENABLE_s1.address
		.TRANSMIT_ENABLE_s1_write                       (mm_interconnect_0_transmit_enable_s1_write),                       //                                    .write
		.TRANSMIT_ENABLE_s1_readdata                    (mm_interconnect_0_transmit_enable_s1_readdata),                    //                                    .readdata
		.TRANSMIT_ENABLE_s1_writedata                   (mm_interconnect_0_transmit_enable_s1_writedata),                   //                                    .writedata
		.TRANSMIT_ENABLE_s1_chipselect                  (mm_interconnect_0_transmit_enable_s1_chipselect),                  //                                    .chipselect
		.TRANSMIT_LOAD_s1_address                       (mm_interconnect_0_transmit_load_s1_address),                       //                    TRANSMIT_LOAD_s1.address
		.TRANSMIT_LOAD_s1_write                         (mm_interconnect_0_transmit_load_s1_write),                         //                                    .write
		.TRANSMIT_LOAD_s1_readdata                      (mm_interconnect_0_transmit_load_s1_readdata),                      //                                    .readdata
		.TRANSMIT_LOAD_s1_writedata                     (mm_interconnect_0_transmit_load_s1_writedata),                     //                                    .writedata
		.TRANSMIT_LOAD_s1_chipselect                    (mm_interconnect_0_transmit_load_s1_chipselect),                    //                                    .chipselect
		.TRANSMIT_PARALLEL_FROM_PROCESSOR_s1_address    (mm_interconnect_0_transmit_parallel_from_processor_s1_address),    // TRANSMIT_PARALLEL_FROM_PROCESSOR_s1.address
		.TRANSMIT_PARALLEL_FROM_PROCESSOR_s1_write      (mm_interconnect_0_transmit_parallel_from_processor_s1_write),      //                                    .write
		.TRANSMIT_PARALLEL_FROM_PROCESSOR_s1_readdata   (mm_interconnect_0_transmit_parallel_from_processor_s1_readdata),   //                                    .readdata
		.TRANSMIT_PARALLEL_FROM_PROCESSOR_s1_writedata  (mm_interconnect_0_transmit_parallel_from_processor_s1_writedata),  //                                    .writedata
		.TRANSMIT_PARALLEL_FROM_PROCESSOR_s1_chipselect (mm_interconnect_0_transmit_parallel_from_processor_s1_chipselect)  //                                    .chipselect
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule

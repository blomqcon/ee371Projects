// lab5CPU.v

// Generated using ACDS version 15.1 189

`timescale 1 ps / 1 ps
module lab5CPU (
		input  wire        alien_shoot_external_connection_export,              //              alien_shoot_external_connection.export
		input  wire [2:0]  alien_x_external_connection_export,                  //                  alien_x_external_connection.export
		input  wire [1:0]  alien_y_external_connection_export,                  //                  alien_y_external_connection.export
		input  wire        character_recieved_input_external_connection_export, // character_recieved_input_external_connection.export
		input  wire        character_sent_input_external_connection_export,     //     character_sent_input_external_connection.export
		input  wire        clk_clk,                                             //                                          clk.clk
		input  wire [31:0] game_time_external_connection_export,                //                game_time_external_connection.export
		input  wire        gun_left_external_connection_export,                 //                 gun_left_external_connection.export
		input  wire        gun_right_external_connection_export,                //                gun_right_external_connection.export
		input  wire [1:0]  gun_shoot_external_connection_export,                //                gun_shoot_external_connection.export
		output wire [7:0]  led_output_external_connection_export,               //               led_output_external_connection.export
		output wire        load_output_external_connection_export,              //              load_output_external_connection.export
		input  wire [7:0]  parallel_input_external_connection_export,           //           parallel_input_external_connection.export
		output wire [7:0]  parallel_output_external_connection_export,          //          parallel_output_external_connection.export
		input  wire [15:0] random_number_external_connection_export,            //            random_number_external_connection.export
		input  wire        reset_reset_n,                                       //                                        reset.reset_n
		output wire [10:0] sram_address_external_connection_export,             //             sram_address_external_connection.export
		inout  wire [7:0]  sram_data_external_connection_export,                //                sram_data_external_connection.export
		output wire        sram_enable_read_external_connection_export,         //         sram_enable_read_external_connection.export
		output wire        sram_enable_write_external_connection_export,        //        sram_enable_write_external_connection.export
		output wire        transmit_enable_output_external_connection_export    //   transmit_enable_output_external_connection.export
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [14:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [14:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;          // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;       // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;       // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;           // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;              // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;        // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;             // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;         // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_mem_s1_chipselect;                // mm_interconnect_0:onchip_mem_s1_chipselect -> onchip_mem:chipselect
	wire  [31:0] mm_interconnect_0_onchip_mem_s1_readdata;                  // onchip_mem:readdata -> mm_interconnect_0:onchip_mem_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_mem_s1_address;                   // mm_interconnect_0:onchip_mem_s1_address -> onchip_mem:address
	wire   [3:0] mm_interconnect_0_onchip_mem_s1_byteenable;                // mm_interconnect_0:onchip_mem_s1_byteenable -> onchip_mem:byteenable
	wire         mm_interconnect_0_onchip_mem_s1_write;                     // mm_interconnect_0:onchip_mem_s1_write -> onchip_mem:write
	wire  [31:0] mm_interconnect_0_onchip_mem_s1_writedata;                 // mm_interconnect_0:onchip_mem_s1_writedata -> onchip_mem:writedata
	wire         mm_interconnect_0_onchip_mem_s1_clken;                     // mm_interconnect_0:onchip_mem_s1_clken -> onchip_mem:clken
	wire  [31:0] mm_interconnect_0_parallel_input_s1_readdata;              // parallel_input:readdata -> mm_interconnect_0:parallel_input_s1_readdata
	wire   [1:0] mm_interconnect_0_parallel_input_s1_address;               // mm_interconnect_0:parallel_input_s1_address -> parallel_input:address
	wire         mm_interconnect_0_character_recieved_input_s1_chipselect;  // mm_interconnect_0:character_recieved_input_s1_chipselect -> character_recieved_input:chipselect
	wire  [31:0] mm_interconnect_0_character_recieved_input_s1_readdata;    // character_recieved_input:readdata -> mm_interconnect_0:character_recieved_input_s1_readdata
	wire   [1:0] mm_interconnect_0_character_recieved_input_s1_address;     // mm_interconnect_0:character_recieved_input_s1_address -> character_recieved_input:address
	wire         mm_interconnect_0_character_recieved_input_s1_write;       // mm_interconnect_0:character_recieved_input_s1_write -> character_recieved_input:write_n
	wire  [31:0] mm_interconnect_0_character_recieved_input_s1_writedata;   // mm_interconnect_0:character_recieved_input_s1_writedata -> character_recieved_input:writedata
	wire         mm_interconnect_0_led_output_s1_chipselect;                // mm_interconnect_0:led_output_s1_chipselect -> led_output:chipselect
	wire  [31:0] mm_interconnect_0_led_output_s1_readdata;                  // led_output:readdata -> mm_interconnect_0:led_output_s1_readdata
	wire   [1:0] mm_interconnect_0_led_output_s1_address;                   // mm_interconnect_0:led_output_s1_address -> led_output:address
	wire         mm_interconnect_0_led_output_s1_write;                     // mm_interconnect_0:led_output_s1_write -> led_output:write_n
	wire  [31:0] mm_interconnect_0_led_output_s1_writedata;                 // mm_interconnect_0:led_output_s1_writedata -> led_output:writedata
	wire         mm_interconnect_0_parallel_output_s1_chipselect;           // mm_interconnect_0:parallel_output_s1_chipselect -> parallel_output:chipselect
	wire  [31:0] mm_interconnect_0_parallel_output_s1_readdata;             // parallel_output:readdata -> mm_interconnect_0:parallel_output_s1_readdata
	wire   [1:0] mm_interconnect_0_parallel_output_s1_address;              // mm_interconnect_0:parallel_output_s1_address -> parallel_output:address
	wire         mm_interconnect_0_parallel_output_s1_write;                // mm_interconnect_0:parallel_output_s1_write -> parallel_output:write_n
	wire  [31:0] mm_interconnect_0_parallel_output_s1_writedata;            // mm_interconnect_0:parallel_output_s1_writedata -> parallel_output:writedata
	wire         mm_interconnect_0_load_output_s1_chipselect;               // mm_interconnect_0:load_output_s1_chipselect -> load_output:chipselect
	wire  [31:0] mm_interconnect_0_load_output_s1_readdata;                 // load_output:readdata -> mm_interconnect_0:load_output_s1_readdata
	wire   [1:0] mm_interconnect_0_load_output_s1_address;                  // mm_interconnect_0:load_output_s1_address -> load_output:address
	wire         mm_interconnect_0_load_output_s1_write;                    // mm_interconnect_0:load_output_s1_write -> load_output:write_n
	wire  [31:0] mm_interconnect_0_load_output_s1_writedata;                // mm_interconnect_0:load_output_s1_writedata -> load_output:writedata
	wire         mm_interconnect_0_character_sent_input_s1_chipselect;      // mm_interconnect_0:character_sent_input_s1_chipselect -> character_sent_input:chipselect
	wire  [31:0] mm_interconnect_0_character_sent_input_s1_readdata;        // character_sent_input:readdata -> mm_interconnect_0:character_sent_input_s1_readdata
	wire   [1:0] mm_interconnect_0_character_sent_input_s1_address;         // mm_interconnect_0:character_sent_input_s1_address -> character_sent_input:address
	wire         mm_interconnect_0_character_sent_input_s1_write;           // mm_interconnect_0:character_sent_input_s1_write -> character_sent_input:write_n
	wire  [31:0] mm_interconnect_0_character_sent_input_s1_writedata;       // mm_interconnect_0:character_sent_input_s1_writedata -> character_sent_input:writedata
	wire         mm_interconnect_0_transmit_enable_output_s1_chipselect;    // mm_interconnect_0:transmit_enable_output_s1_chipselect -> transmit_enable_output:chipselect
	wire  [31:0] mm_interconnect_0_transmit_enable_output_s1_readdata;      // transmit_enable_output:readdata -> mm_interconnect_0:transmit_enable_output_s1_readdata
	wire   [1:0] mm_interconnect_0_transmit_enable_output_s1_address;       // mm_interconnect_0:transmit_enable_output_s1_address -> transmit_enable_output:address
	wire         mm_interconnect_0_transmit_enable_output_s1_write;         // mm_interconnect_0:transmit_enable_output_s1_write -> transmit_enable_output:write_n
	wire  [31:0] mm_interconnect_0_transmit_enable_output_s1_writedata;     // mm_interconnect_0:transmit_enable_output_s1_writedata -> transmit_enable_output:writedata
	wire         mm_interconnect_0_sram_data_s1_chipselect;                 // mm_interconnect_0:sram_data_s1_chipselect -> sram_data:chipselect
	wire  [31:0] mm_interconnect_0_sram_data_s1_readdata;                   // sram_data:readdata -> mm_interconnect_0:sram_data_s1_readdata
	wire   [1:0] mm_interconnect_0_sram_data_s1_address;                    // mm_interconnect_0:sram_data_s1_address -> sram_data:address
	wire         mm_interconnect_0_sram_data_s1_write;                      // mm_interconnect_0:sram_data_s1_write -> sram_data:write_n
	wire  [31:0] mm_interconnect_0_sram_data_s1_writedata;                  // mm_interconnect_0:sram_data_s1_writedata -> sram_data:writedata
	wire         mm_interconnect_0_sram_enable_write_s1_chipselect;         // mm_interconnect_0:sram_enable_write_s1_chipselect -> sram_enable_write:chipselect
	wire  [31:0] mm_interconnect_0_sram_enable_write_s1_readdata;           // sram_enable_write:readdata -> mm_interconnect_0:sram_enable_write_s1_readdata
	wire   [1:0] mm_interconnect_0_sram_enable_write_s1_address;            // mm_interconnect_0:sram_enable_write_s1_address -> sram_enable_write:address
	wire         mm_interconnect_0_sram_enable_write_s1_write;              // mm_interconnect_0:sram_enable_write_s1_write -> sram_enable_write:write_n
	wire  [31:0] mm_interconnect_0_sram_enable_write_s1_writedata;          // mm_interconnect_0:sram_enable_write_s1_writedata -> sram_enable_write:writedata
	wire         mm_interconnect_0_sram_enable_read_s1_chipselect;          // mm_interconnect_0:sram_enable_read_s1_chipselect -> sram_enable_read:chipselect
	wire  [31:0] mm_interconnect_0_sram_enable_read_s1_readdata;            // sram_enable_read:readdata -> mm_interconnect_0:sram_enable_read_s1_readdata
	wire   [1:0] mm_interconnect_0_sram_enable_read_s1_address;             // mm_interconnect_0:sram_enable_read_s1_address -> sram_enable_read:address
	wire         mm_interconnect_0_sram_enable_read_s1_write;               // mm_interconnect_0:sram_enable_read_s1_write -> sram_enable_read:write_n
	wire  [31:0] mm_interconnect_0_sram_enable_read_s1_writedata;           // mm_interconnect_0:sram_enable_read_s1_writedata -> sram_enable_read:writedata
	wire         mm_interconnect_0_sram_address_s1_chipselect;              // mm_interconnect_0:sram_address_s1_chipselect -> sram_address:chipselect
	wire  [31:0] mm_interconnect_0_sram_address_s1_readdata;                // sram_address:readdata -> mm_interconnect_0:sram_address_s1_readdata
	wire   [1:0] mm_interconnect_0_sram_address_s1_address;                 // mm_interconnect_0:sram_address_s1_address -> sram_address:address
	wire         mm_interconnect_0_sram_address_s1_write;                   // mm_interconnect_0:sram_address_s1_write -> sram_address:write_n
	wire  [31:0] mm_interconnect_0_sram_address_s1_writedata;               // mm_interconnect_0:sram_address_s1_writedata -> sram_address:writedata
	wire         mm_interconnect_0_gun_left_s1_chipselect;                  // mm_interconnect_0:gun_left_s1_chipselect -> gun_left:chipselect
	wire  [31:0] mm_interconnect_0_gun_left_s1_readdata;                    // gun_left:readdata -> mm_interconnect_0:gun_left_s1_readdata
	wire   [1:0] mm_interconnect_0_gun_left_s1_address;                     // mm_interconnect_0:gun_left_s1_address -> gun_left:address
	wire         mm_interconnect_0_gun_left_s1_write;                       // mm_interconnect_0:gun_left_s1_write -> gun_left:write_n
	wire  [31:0] mm_interconnect_0_gun_left_s1_writedata;                   // mm_interconnect_0:gun_left_s1_writedata -> gun_left:writedata
	wire         mm_interconnect_0_gun_right_s1_chipselect;                 // mm_interconnect_0:gun_right_s1_chipselect -> gun_right:chipselect
	wire  [31:0] mm_interconnect_0_gun_right_s1_readdata;                   // gun_right:readdata -> mm_interconnect_0:gun_right_s1_readdata
	wire   [1:0] mm_interconnect_0_gun_right_s1_address;                    // mm_interconnect_0:gun_right_s1_address -> gun_right:address
	wire         mm_interconnect_0_gun_right_s1_write;                      // mm_interconnect_0:gun_right_s1_write -> gun_right:write_n
	wire  [31:0] mm_interconnect_0_gun_right_s1_writedata;                  // mm_interconnect_0:gun_right_s1_writedata -> gun_right:writedata
	wire         mm_interconnect_0_gun_shoot_s1_chipselect;                 // mm_interconnect_0:gun_shoot_s1_chipselect -> gun_shoot:chipselect
	wire  [31:0] mm_interconnect_0_gun_shoot_s1_readdata;                   // gun_shoot:readdata -> mm_interconnect_0:gun_shoot_s1_readdata
	wire   [1:0] mm_interconnect_0_gun_shoot_s1_address;                    // mm_interconnect_0:gun_shoot_s1_address -> gun_shoot:address
	wire         mm_interconnect_0_gun_shoot_s1_write;                      // mm_interconnect_0:gun_shoot_s1_write -> gun_shoot:write_n
	wire  [31:0] mm_interconnect_0_gun_shoot_s1_writedata;                  // mm_interconnect_0:gun_shoot_s1_writedata -> gun_shoot:writedata
	wire  [31:0] mm_interconnect_0_alien_x_s1_readdata;                     // alien_x:readdata -> mm_interconnect_0:alien_x_s1_readdata
	wire   [1:0] mm_interconnect_0_alien_x_s1_address;                      // mm_interconnect_0:alien_x_s1_address -> alien_x:address
	wire  [31:0] mm_interconnect_0_alien_y_s1_readdata;                     // alien_y:readdata -> mm_interconnect_0:alien_y_s1_readdata
	wire   [1:0] mm_interconnect_0_alien_y_s1_address;                      // mm_interconnect_0:alien_y_s1_address -> alien_y:address
	wire  [31:0] mm_interconnect_0_alien_shoot_s1_readdata;                 // alien_shoot:readdata -> mm_interconnect_0:alien_shoot_s1_readdata
	wire   [1:0] mm_interconnect_0_alien_shoot_s1_address;                  // mm_interconnect_0:alien_shoot_s1_address -> alien_shoot:address
	wire  [31:0] mm_interconnect_0_random_number_s1_readdata;               // random_number:readdata -> mm_interconnect_0:random_number_s1_readdata
	wire   [1:0] mm_interconnect_0_random_number_s1_address;                // mm_interconnect_0:random_number_s1_address -> random_number:address
	wire  [31:0] mm_interconnect_0_game_time_s1_readdata;                   // game_time:readdata -> mm_interconnect_0:game_time_s1_readdata
	wire   [1:0] mm_interconnect_0_game_time_s1_address;                    // mm_interconnect_0:game_time_s1_address -> game_time:address
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // gun_left:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // character_recieved_input:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // character_sent_input:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // gun_right:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                  // gun_shoot:irq -> irq_mapper:receiver5_irq
	wire  [31:0] cpu_d_irq_irq;                                             // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [alien_shoot:reset_n, alien_x:reset_n, alien_y:reset_n, character_recieved_input:reset_n, character_sent_input:reset_n, cpu:reset_n, game_time:reset_n, gun_left:reset_n, gun_right:reset_n, gun_shoot:reset_n, irq_mapper:reset, jtag_uart:rst_n, led_output:reset_n, load_output:reset_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_mem:reset, parallel_input:reset_n, parallel_output:reset_n, random_number:reset_n, rst_translator:in_reset, sram_address:reset_n, sram_data:reset_n, sram_enable_read:reset_n, sram_enable_write:reset_n, transmit_enable_output:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, onchip_mem:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                         // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	lab5CPU_alien_shoot alien_shoot (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_alien_shoot_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_alien_shoot_s1_readdata), //                    .readdata
		.in_port  (alien_shoot_external_connection_export)     // external_connection.export
	);

	lab5CPU_alien_x alien_x (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_alien_x_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_alien_x_s1_readdata), //                    .readdata
		.in_port  (alien_x_external_connection_export)     // external_connection.export
	);

	lab5CPU_alien_y alien_y (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_alien_y_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_alien_y_s1_readdata), //                    .readdata
		.in_port  (alien_y_external_connection_export)     // external_connection.export
	);

	lab5CPU_character_recieved_input character_recieved_input (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                          //               reset.reset_n
		.address    (mm_interconnect_0_character_recieved_input_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_character_recieved_input_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_character_recieved_input_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_character_recieved_input_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_character_recieved_input_s1_readdata),   //                    .readdata
		.in_port    (character_recieved_input_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                                  //                 irq.irq
	);

	lab5CPU_character_recieved_input character_sent_input (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (mm_interconnect_0_character_sent_input_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_character_sent_input_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_character_sent_input_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_character_sent_input_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_character_sent_input_s1_readdata),   //                    .readdata
		.in_port    (character_sent_input_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                              //                 irq.irq
	);

	lab5CPU_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	lab5CPU_game_time game_time (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_game_time_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_game_time_s1_readdata), //                    .readdata
		.in_port  (game_time_external_connection_export)     // external_connection.export
	);

	lab5CPU_character_recieved_input gun_left (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_gun_left_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gun_left_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gun_left_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gun_left_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gun_left_s1_readdata),   //                    .readdata
		.in_port    (gun_left_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                  //                 irq.irq
	);

	lab5CPU_character_recieved_input gun_right (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_gun_right_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gun_right_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gun_right_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gun_right_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gun_right_s1_readdata),   //                    .readdata
		.in_port    (gun_right_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                   //                 irq.irq
	);

	lab5CPU_gun_shoot gun_shoot (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_gun_shoot_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gun_shoot_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gun_shoot_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gun_shoot_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gun_shoot_s1_readdata),   //                    .readdata
		.in_port    (gun_shoot_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                   //                 irq.irq
	);

	lab5CPU_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	lab5CPU_led_output led_output (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_led_output_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_output_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_output_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_output_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_output_s1_readdata),   //                    .readdata
		.out_port   (led_output_external_connection_export)       // external_connection.export
	);

	lab5CPU_load_output load_output (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_load_output_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_load_output_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_load_output_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_load_output_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_load_output_s1_readdata),   //                    .readdata
		.out_port   (load_output_external_connection_export)       // external_connection.export
	);

	lab5CPU_onchip_mem onchip_mem (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	lab5CPU_parallel_input parallel_input (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_parallel_input_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_parallel_input_s1_readdata), //                    .readdata
		.in_port  (parallel_input_external_connection_export)     // external_connection.export
	);

	lab5CPU_led_output parallel_output (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_parallel_output_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_parallel_output_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_parallel_output_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_parallel_output_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_parallel_output_s1_readdata),   //                    .readdata
		.out_port   (parallel_output_external_connection_export)       // external_connection.export
	);

	lab5CPU_random_number random_number (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_random_number_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_random_number_s1_readdata), //                    .readdata
		.in_port  (random_number_external_connection_export)     // external_connection.export
	);

	lab5CPU_sram_address sram_address (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_sram_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sram_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sram_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sram_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sram_address_s1_readdata),   //                    .readdata
		.out_port   (sram_address_external_connection_export)       // external_connection.export
	);

	lab5CPU_sram_data sram_data (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_sram_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sram_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sram_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sram_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sram_data_s1_readdata),   //                    .readdata
		.bidir_port (sram_data_external_connection_export)       // external_connection.export
	);

	lab5CPU_load_output sram_enable_read (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_sram_enable_read_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sram_enable_read_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sram_enable_read_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sram_enable_read_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sram_enable_read_s1_readdata),   //                    .readdata
		.out_port   (sram_enable_read_external_connection_export)       // external_connection.export
	);

	lab5CPU_load_output sram_enable_write (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_sram_enable_write_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sram_enable_write_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sram_enable_write_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sram_enable_write_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sram_enable_write_s1_readdata),   //                    .readdata
		.out_port   (sram_enable_write_external_connection_export)       // external_connection.export
	);

	lab5CPU_load_output transmit_enable_output (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (mm_interconnect_0_transmit_enable_output_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_transmit_enable_output_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_transmit_enable_output_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_transmit_enable_output_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_transmit_enable_output_s1_readdata),   //                    .readdata
		.out_port   (transmit_enable_output_external_connection_export)       // external_connection.export
	);

	lab5CPU_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                           (clk_clk),                                                   //                         clk_0_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                   cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                  .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                  .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                  .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                  .readdata
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                  .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                  .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                  .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //            cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                  .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                  .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                  .readdata
		.alien_shoot_s1_address                  (mm_interconnect_0_alien_shoot_s1_address),                  //                    alien_shoot_s1.address
		.alien_shoot_s1_readdata                 (mm_interconnect_0_alien_shoot_s1_readdata),                 //                                  .readdata
		.alien_x_s1_address                      (mm_interconnect_0_alien_x_s1_address),                      //                        alien_x_s1.address
		.alien_x_s1_readdata                     (mm_interconnect_0_alien_x_s1_readdata),                     //                                  .readdata
		.alien_y_s1_address                      (mm_interconnect_0_alien_y_s1_address),                      //                        alien_y_s1.address
		.alien_y_s1_readdata                     (mm_interconnect_0_alien_y_s1_readdata),                     //                                  .readdata
		.character_recieved_input_s1_address     (mm_interconnect_0_character_recieved_input_s1_address),     //       character_recieved_input_s1.address
		.character_recieved_input_s1_write       (mm_interconnect_0_character_recieved_input_s1_write),       //                                  .write
		.character_recieved_input_s1_readdata    (mm_interconnect_0_character_recieved_input_s1_readdata),    //                                  .readdata
		.character_recieved_input_s1_writedata   (mm_interconnect_0_character_recieved_input_s1_writedata),   //                                  .writedata
		.character_recieved_input_s1_chipselect  (mm_interconnect_0_character_recieved_input_s1_chipselect),  //                                  .chipselect
		.character_sent_input_s1_address         (mm_interconnect_0_character_sent_input_s1_address),         //           character_sent_input_s1.address
		.character_sent_input_s1_write           (mm_interconnect_0_character_sent_input_s1_write),           //                                  .write
		.character_sent_input_s1_readdata        (mm_interconnect_0_character_sent_input_s1_readdata),        //                                  .readdata
		.character_sent_input_s1_writedata       (mm_interconnect_0_character_sent_input_s1_writedata),       //                                  .writedata
		.character_sent_input_s1_chipselect      (mm_interconnect_0_character_sent_input_s1_chipselect),      //                                  .chipselect
		.cpu_jtag_debug_module_address           (mm_interconnect_0_cpu_jtag_debug_module_address),           //             cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write             (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                  .write
		.cpu_jtag_debug_module_read              (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                  .read
		.cpu_jtag_debug_module_readdata          (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                  .readdata
		.cpu_jtag_debug_module_writedata         (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                  .writedata
		.cpu_jtag_debug_module_byteenable        (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                  .byteenable
		.cpu_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                  .waitrequest
		.cpu_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                  .debugaccess
		.game_time_s1_address                    (mm_interconnect_0_game_time_s1_address),                    //                      game_time_s1.address
		.game_time_s1_readdata                   (mm_interconnect_0_game_time_s1_readdata),                   //                                  .readdata
		.gun_left_s1_address                     (mm_interconnect_0_gun_left_s1_address),                     //                       gun_left_s1.address
		.gun_left_s1_write                       (mm_interconnect_0_gun_left_s1_write),                       //                                  .write
		.gun_left_s1_readdata                    (mm_interconnect_0_gun_left_s1_readdata),                    //                                  .readdata
		.gun_left_s1_writedata                   (mm_interconnect_0_gun_left_s1_writedata),                   //                                  .writedata
		.gun_left_s1_chipselect                  (mm_interconnect_0_gun_left_s1_chipselect),                  //                                  .chipselect
		.gun_right_s1_address                    (mm_interconnect_0_gun_right_s1_address),                    //                      gun_right_s1.address
		.gun_right_s1_write                      (mm_interconnect_0_gun_right_s1_write),                      //                                  .write
		.gun_right_s1_readdata                   (mm_interconnect_0_gun_right_s1_readdata),                   //                                  .readdata
		.gun_right_s1_writedata                  (mm_interconnect_0_gun_right_s1_writedata),                  //                                  .writedata
		.gun_right_s1_chipselect                 (mm_interconnect_0_gun_right_s1_chipselect),                 //                                  .chipselect
		.gun_shoot_s1_address                    (mm_interconnect_0_gun_shoot_s1_address),                    //                      gun_shoot_s1.address
		.gun_shoot_s1_write                      (mm_interconnect_0_gun_shoot_s1_write),                      //                                  .write
		.gun_shoot_s1_readdata                   (mm_interconnect_0_gun_shoot_s1_readdata),                   //                                  .readdata
		.gun_shoot_s1_writedata                  (mm_interconnect_0_gun_shoot_s1_writedata),                  //                                  .writedata
		.gun_shoot_s1_chipselect                 (mm_interconnect_0_gun_shoot_s1_chipselect),                 //                                  .chipselect
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.led_output_s1_address                   (mm_interconnect_0_led_output_s1_address),                   //                     led_output_s1.address
		.led_output_s1_write                     (mm_interconnect_0_led_output_s1_write),                     //                                  .write
		.led_output_s1_readdata                  (mm_interconnect_0_led_output_s1_readdata),                  //                                  .readdata
		.led_output_s1_writedata                 (mm_interconnect_0_led_output_s1_writedata),                 //                                  .writedata
		.led_output_s1_chipselect                (mm_interconnect_0_led_output_s1_chipselect),                //                                  .chipselect
		.load_output_s1_address                  (mm_interconnect_0_load_output_s1_address),                  //                    load_output_s1.address
		.load_output_s1_write                    (mm_interconnect_0_load_output_s1_write),                    //                                  .write
		.load_output_s1_readdata                 (mm_interconnect_0_load_output_s1_readdata),                 //                                  .readdata
		.load_output_s1_writedata                (mm_interconnect_0_load_output_s1_writedata),                //                                  .writedata
		.load_output_s1_chipselect               (mm_interconnect_0_load_output_s1_chipselect),               //                                  .chipselect
		.onchip_mem_s1_address                   (mm_interconnect_0_onchip_mem_s1_address),                   //                     onchip_mem_s1.address
		.onchip_mem_s1_write                     (mm_interconnect_0_onchip_mem_s1_write),                     //                                  .write
		.onchip_mem_s1_readdata                  (mm_interconnect_0_onchip_mem_s1_readdata),                  //                                  .readdata
		.onchip_mem_s1_writedata                 (mm_interconnect_0_onchip_mem_s1_writedata),                 //                                  .writedata
		.onchip_mem_s1_byteenable                (mm_interconnect_0_onchip_mem_s1_byteenable),                //                                  .byteenable
		.onchip_mem_s1_chipselect                (mm_interconnect_0_onchip_mem_s1_chipselect),                //                                  .chipselect
		.onchip_mem_s1_clken                     (mm_interconnect_0_onchip_mem_s1_clken),                     //                                  .clken
		.parallel_input_s1_address               (mm_interconnect_0_parallel_input_s1_address),               //                 parallel_input_s1.address
		.parallel_input_s1_readdata              (mm_interconnect_0_parallel_input_s1_readdata),              //                                  .readdata
		.parallel_output_s1_address              (mm_interconnect_0_parallel_output_s1_address),              //                parallel_output_s1.address
		.parallel_output_s1_write                (mm_interconnect_0_parallel_output_s1_write),                //                                  .write
		.parallel_output_s1_readdata             (mm_interconnect_0_parallel_output_s1_readdata),             //                                  .readdata
		.parallel_output_s1_writedata            (mm_interconnect_0_parallel_output_s1_writedata),            //                                  .writedata
		.parallel_output_s1_chipselect           (mm_interconnect_0_parallel_output_s1_chipselect),           //                                  .chipselect
		.random_number_s1_address                (mm_interconnect_0_random_number_s1_address),                //                  random_number_s1.address
		.random_number_s1_readdata               (mm_interconnect_0_random_number_s1_readdata),               //                                  .readdata
		.sram_address_s1_address                 (mm_interconnect_0_sram_address_s1_address),                 //                   sram_address_s1.address
		.sram_address_s1_write                   (mm_interconnect_0_sram_address_s1_write),                   //                                  .write
		.sram_address_s1_readdata                (mm_interconnect_0_sram_address_s1_readdata),                //                                  .readdata
		.sram_address_s1_writedata               (mm_interconnect_0_sram_address_s1_writedata),               //                                  .writedata
		.sram_address_s1_chipselect              (mm_interconnect_0_sram_address_s1_chipselect),              //                                  .chipselect
		.sram_data_s1_address                    (mm_interconnect_0_sram_data_s1_address),                    //                      sram_data_s1.address
		.sram_data_s1_write                      (mm_interconnect_0_sram_data_s1_write),                      //                                  .write
		.sram_data_s1_readdata                   (mm_interconnect_0_sram_data_s1_readdata),                   //                                  .readdata
		.sram_data_s1_writedata                  (mm_interconnect_0_sram_data_s1_writedata),                  //                                  .writedata
		.sram_data_s1_chipselect                 (mm_interconnect_0_sram_data_s1_chipselect),                 //                                  .chipselect
		.sram_enable_read_s1_address             (mm_interconnect_0_sram_enable_read_s1_address),             //               sram_enable_read_s1.address
		.sram_enable_read_s1_write               (mm_interconnect_0_sram_enable_read_s1_write),               //                                  .write
		.sram_enable_read_s1_readdata            (mm_interconnect_0_sram_enable_read_s1_readdata),            //                                  .readdata
		.sram_enable_read_s1_writedata           (mm_interconnect_0_sram_enable_read_s1_writedata),           //                                  .writedata
		.sram_enable_read_s1_chipselect          (mm_interconnect_0_sram_enable_read_s1_chipselect),          //                                  .chipselect
		.sram_enable_write_s1_address            (mm_interconnect_0_sram_enable_write_s1_address),            //              sram_enable_write_s1.address
		.sram_enable_write_s1_write              (mm_interconnect_0_sram_enable_write_s1_write),              //                                  .write
		.sram_enable_write_s1_readdata           (mm_interconnect_0_sram_enable_write_s1_readdata),           //                                  .readdata
		.sram_enable_write_s1_writedata          (mm_interconnect_0_sram_enable_write_s1_writedata),          //                                  .writedata
		.sram_enable_write_s1_chipselect         (mm_interconnect_0_sram_enable_write_s1_chipselect),         //                                  .chipselect
		.transmit_enable_output_s1_address       (mm_interconnect_0_transmit_enable_output_s1_address),       //         transmit_enable_output_s1.address
		.transmit_enable_output_s1_write         (mm_interconnect_0_transmit_enable_output_s1_write),         //                                  .write
		.transmit_enable_output_s1_readdata      (mm_interconnect_0_transmit_enable_output_s1_readdata),      //                                  .readdata
		.transmit_enable_output_s1_writedata     (mm_interconnect_0_transmit_enable_output_s1_writedata),     //                                  .writedata
		.transmit_enable_output_s1_chipselect    (mm_interconnect_0_transmit_enable_output_s1_chipselect)     //                                  .chipselect
	);

	lab5CPU_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
